------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity trigger is
    generic(
        g_NUM_OF_OHs : integer := 1
    );
    port(
        -- reset
        reset_i             : in  std_logic;
        
        -- TTC
        ttc_clk_i           : in  t_ttc_clks;
        ttc_cmds_i          : in  t_ttc_cmds;

        -- Sbit cluster inputs
        sbit_clusters_i     : in t_oh_sbits_arr(g_NUM_OF_OHs - 1 downto 0);
        sbit_link_status_i  : in t_oh_sbit_links_arr(g_NUM_OF_OHs - 1 downto 0);

        -- Outputs
        trig_led_o          : out std_logic;

        -- IPbus
        ipb_reset_i         : in  std_logic;
        ipb_clk_i           : in  std_logic;
        ipb_miso_o          : out ipb_rbus;
        ipb_mosi_i          : in  ipb_wbus
    );
end trigger;

architecture trigger_arch of trigger is
    
    signal reset_global         : std_logic;
    signal reset_local          : std_logic;
    signal reset                : std_logic;
    signal reset_cnt            : std_logic;
    
    signal oh_mask              : std_logic_vector(23 downto 0) := (others => '0');
    signal oh_triggers          : std_logic_vector(g_NUM_OF_OHs - 1 downto 0) := (others => '0');
    signal or_trigger           : std_logic;
        
    signal sbitmon_reset        : std_logic;
    signal sbitmon_sbits        : t_oh_sbits;
    signal sbitmon_link_select  : std_logic_vector(3 downto 0);
    
    -- counters
    signal or_trigger_rate      : std_logic_vector(31 downto 0); 
    signal or_trigger_cnt       : std_logic_vector(31 downto 0); 
    
    -- OH counters
    signal sbit_overflow_cnt    : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal missed_comma_cnt     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal link_overflow_cnt    : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal link_underflow_cnt   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_word_cnt        : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trigger_rate         : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trigger_cnt          : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal cluster_cnt_rate     : t_std32_array((g_NUM_OF_OHs * 9) - 1 downto 0);
    signal cluster_cnt          : t_std32_array((g_NUM_OF_OHs * 9) - 1 downto 0);
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_TRIGGER_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;

    --== Trigger ==--
    
    or_trigger <= or_reduce(oh_triggers);

    i_or_trigger_rate : entity work.rate_counter
        generic map(
            g_CLK_FREQUENCY => C_TTC_CLK_FREQUENCY_SLV,
            g_COUNTER_WIDTH => 32
        )
        port map(
            clk_i   => ttc_clk_i.clk_40,
            reset_i => reset or reset_cnt,
            en_i    => or_trigger,
            rate_o  => or_trigger_rate
        );

    i_or_trigger_cnt: entity work.counter
        generic map(
            g_COUNTER_WIDTH  => 32,
            g_ALLOW_ROLLOVER => FALSE
        )
        port map(
            ref_clk_i => ttc_clk_i.clk_40,
            reset_i   => reset or reset_cnt,
            en_i      => or_trigger,
            count_o   => or_trigger_cnt
        );
    
    i_led_pulse : entity work.pulse_extend
        generic map(
            DELAY_CNT_LENGTH => C_LED_PULSE_LENGTH_TTC_CLK'length
        )
        port map(
            clk_i          => ttc_clk_i.clk_40,
            rst_i          => reset,
            pulse_length_i => C_LED_PULSE_LENGTH_TTC_CLK,
            pulse_i        => or_trigger,
            pulse_o        => trig_led_o
        );
    
    --== Links ==--
        
    -- TODO: imlpement link synchronization by looking for sync words after each resync and delay the data of all links to match the latest one (use FIFOs for that) 
    g_input_processors:
    for i in 0 to g_NUM_OF_OHs - 1 generate
        
        i_input_processor: entity work.trigger_input_processor
            port map(
                reset_i              => reset,
                reset_cnt_i          => reset_cnt,
                clk_i                => ttc_clk_i.clk_40,
                sbit_clusters_i      => sbit_clusters_i(i),
                link_status_i        => sbit_link_status_i(i),
                masked_i             => oh_mask(i),
                trigger_o            => oh_triggers(i),
                sbit_overflow_cnt_o  => sbit_overflow_cnt(i),
                missed_comma_cnt_o   => missed_comma_cnt(i),
                link_overflow_cnt_o  => link_overflow_cnt(i),
                link_underflow_cnt_o => link_underflow_cnt(i),
                sync_word_cnt_o      => sync_word_cnt(i),
                cluster_cnt_rate_o   => cluster_cnt_rate(((i + 1) * 9) - 1 downto i * 9),
                trigger_rate_o       => trigger_rate(i),
                cluster_cnt_o        => cluster_cnt(((i + 1) * 9) - 1 downto i * 9),
                trigger_cnt_o        => trigger_cnt(i)
            );
        
    end generate;

    --== SBit monitor ==--
    
    i_sbit_monitor : entity work.sbit_monitor
        generic map(
            g_NUM_OF_OHs => g_NUM_OF_OHs
        )
        port map(
            reset_i         => sbitmon_reset,
            ttc_clk_i       => ttc_clk_i,
            link_select_i   => sbitmon_link_select,
            sbit_clusters_i => sbit_clusters_i,
            sbit_trigger_i  => oh_triggers,
            frozen_sbits_o  => sbitmon_sbits
        );
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_TRIGGER_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_TRIGGER_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_TRIGGER_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"000";
    regs_addresses(1)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"001";
    regs_addresses(2)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"002";
    regs_addresses(3)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"010";
    regs_addresses(4)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"011";
    regs_addresses(5)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"080";
    regs_addresses(6)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"081";
    regs_addresses(7)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"082";
    regs_addresses(8)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"083";
    regs_addresses(9)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"084";
    regs_addresses(10)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"085";
    regs_addresses(11)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"086";
    regs_addresses(12)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"087";
    regs_addresses(13)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"088";
    regs_addresses(14)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"089";
    regs_addresses(15)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"100";
    regs_addresses(16)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"101";
    regs_addresses(17)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"110";
    regs_addresses(18)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"111";
    regs_addresses(19)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"112";
    regs_addresses(20)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"113";
    regs_addresses(21)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"114";
    regs_addresses(22)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"115";
    regs_addresses(23)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"116";
    regs_addresses(24)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"117";
    regs_addresses(25)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"118";
    regs_addresses(26)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"120";
    regs_addresses(27)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"121";
    regs_addresses(28)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"122";
    regs_addresses(29)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"123";
    regs_addresses(30)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"124";
    regs_addresses(31)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"125";
    regs_addresses(32)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"126";
    regs_addresses(33)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"127";
    regs_addresses(34)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"128";
    regs_addresses(35)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a0";
    regs_addresses(36)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a1";
    regs_addresses(37)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a3";
    regs_addresses(38)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a4";
    regs_addresses(39)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"1a5";
    regs_addresses(40)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"200";
    regs_addresses(41)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"201";
    regs_addresses(42)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"210";
    regs_addresses(43)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"211";
    regs_addresses(44)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"212";
    regs_addresses(45)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"213";
    regs_addresses(46)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"214";
    regs_addresses(47)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"215";
    regs_addresses(48)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"216";
    regs_addresses(49)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"217";
    regs_addresses(50)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"218";
    regs_addresses(51)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"220";
    regs_addresses(52)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"221";
    regs_addresses(53)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"222";
    regs_addresses(54)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"223";
    regs_addresses(55)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"224";
    regs_addresses(56)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"225";
    regs_addresses(57)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"226";
    regs_addresses(58)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"227";
    regs_addresses(59)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"228";
    regs_addresses(60)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a0";
    regs_addresses(61)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a1";
    regs_addresses(62)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a3";
    regs_addresses(63)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a4";
    regs_addresses(64)(REG_TRIGGER_ADDRESS_MSB downto REG_TRIGGER_ADDRESS_LSB) <= '0' & x"2a5";

    -- Connect read signals
    regs_read_arr(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB) <= oh_mask;
    regs_read_arr(3)(REG_TRIGGER_STATUS_OR_TRIGGER_RATE_MSB downto REG_TRIGGER_STATUS_OR_TRIGGER_RATE_LSB) <= or_trigger_rate;
    regs_read_arr(4)(REG_TRIGGER_STATUS_OR_TRIGGER_CNT_MSB downto REG_TRIGGER_STATUS_OR_TRIGGER_CNT_LSB) <= or_trigger_cnt;
    regs_read_arr(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB) <= sbitmon_link_select;
    regs_read_arr(7)(REG_TRIGGER_SBIT_MONITOR_CLUSTER0_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER0_LSB) <= '0' & sbitmon_sbits(0).size & '0' & sbitmon_sbits(0).address;
    regs_read_arr(8)(REG_TRIGGER_SBIT_MONITOR_CLUSTER1_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER1_LSB) <= '0' & sbitmon_sbits(1).size & '0' & sbitmon_sbits(1).address;
    regs_read_arr(9)(REG_TRIGGER_SBIT_MONITOR_CLUSTER2_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER2_LSB) <= '0' & sbitmon_sbits(2).size & '0' & sbitmon_sbits(2).address;
    regs_read_arr(10)(REG_TRIGGER_SBIT_MONITOR_CLUSTER3_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER3_LSB) <= '0' & sbitmon_sbits(3).size & '0' & sbitmon_sbits(3).address;
    regs_read_arr(11)(REG_TRIGGER_SBIT_MONITOR_CLUSTER4_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER4_LSB) <= '0' & sbitmon_sbits(4).size & '0' & sbitmon_sbits(4).address;
    regs_read_arr(12)(REG_TRIGGER_SBIT_MONITOR_CLUSTER5_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER5_LSB) <= '0' & sbitmon_sbits(5).size & '0' & sbitmon_sbits(5).address;
    regs_read_arr(13)(REG_TRIGGER_SBIT_MONITOR_CLUSTER6_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER6_LSB) <= '0' & sbitmon_sbits(6).size & '0' & sbitmon_sbits(6).address;
    regs_read_arr(14)(REG_TRIGGER_SBIT_MONITOR_CLUSTER7_MSB downto REG_TRIGGER_SBIT_MONITOR_CLUSTER7_LSB) <= '0' & sbitmon_sbits(7).size & '0' & sbitmon_sbits(7).address;
    regs_read_arr(15)(REG_TRIGGER_OH0_TRIGGER_RATE_MSB downto REG_TRIGGER_OH0_TRIGGER_RATE_LSB) <= trigger_rate(0);
    regs_read_arr(16)(REG_TRIGGER_OH0_TRIGGER_CNT_MSB downto REG_TRIGGER_OH0_TRIGGER_CNT_LSB) <= trigger_cnt(0);
    regs_read_arr(17)(REG_TRIGGER_OH0_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 0);
    regs_read_arr(18)(REG_TRIGGER_OH0_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 1);
    regs_read_arr(19)(REG_TRIGGER_OH0_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 2);
    regs_read_arr(20)(REG_TRIGGER_OH0_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 3);
    regs_read_arr(21)(REG_TRIGGER_OH0_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 4);
    regs_read_arr(22)(REG_TRIGGER_OH0_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 5);
    regs_read_arr(23)(REG_TRIGGER_OH0_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 6);
    regs_read_arr(24)(REG_TRIGGER_OH0_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 7);
    regs_read_arr(25)(REG_TRIGGER_OH0_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(0 * 9 + 8);
    regs_read_arr(26)(REG_TRIGGER_OH0_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(0 * 9 + 0);
    regs_read_arr(27)(REG_TRIGGER_OH0_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(0 * 9 + 1);
    regs_read_arr(28)(REG_TRIGGER_OH0_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(0 * 9 + 2);
    regs_read_arr(29)(REG_TRIGGER_OH0_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(0 * 9 + 3);
    regs_read_arr(30)(REG_TRIGGER_OH0_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(0 * 9 + 4);
    regs_read_arr(31)(REG_TRIGGER_OH0_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(0 * 9 + 5);
    regs_read_arr(32)(REG_TRIGGER_OH0_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(0 * 9 + 6);
    regs_read_arr(33)(REG_TRIGGER_OH0_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(0 * 9 + 7);
    regs_read_arr(34)(REG_TRIGGER_OH0_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH0_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(0 * 9 + 8);
    regs_read_arr(35)(REG_TRIGGER_OH0_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(0)(15 downto 0);
    regs_read_arr(35)(REG_TRIGGER_OH0_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(0)(31 downto 16);
    regs_read_arr(36)(REG_TRIGGER_OH0_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH0_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(0)(15 downto 0);
    regs_read_arr(36)(REG_TRIGGER_OH0_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH0_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(0)(31 downto 16);
    regs_read_arr(37)(REG_TRIGGER_OH0_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(0)(15 downto 0);
    regs_read_arr(37)(REG_TRIGGER_OH0_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(0)(31 downto 16);
    regs_read_arr(38)(REG_TRIGGER_OH0_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(0)(15 downto 0);
    regs_read_arr(38)(REG_TRIGGER_OH0_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH0_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(0)(31 downto 16);
    regs_read_arr(39)(REG_TRIGGER_OH0_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH0_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(0)(15 downto 0);
    regs_read_arr(39)(REG_TRIGGER_OH0_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH0_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(0)(31 downto 16);
    regs_read_arr(40)(REG_TRIGGER_OH1_TRIGGER_RATE_MSB downto REG_TRIGGER_OH1_TRIGGER_RATE_LSB) <= trigger_rate(1);
    regs_read_arr(41)(REG_TRIGGER_OH1_TRIGGER_CNT_MSB downto REG_TRIGGER_OH1_TRIGGER_CNT_LSB) <= trigger_cnt(1);
    regs_read_arr(42)(REG_TRIGGER_OH1_CLUSTER_SIZE_0_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_0_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 0);
    regs_read_arr(43)(REG_TRIGGER_OH1_CLUSTER_SIZE_1_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_1_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 1);
    regs_read_arr(44)(REG_TRIGGER_OH1_CLUSTER_SIZE_2_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_2_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 2);
    regs_read_arr(45)(REG_TRIGGER_OH1_CLUSTER_SIZE_3_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_3_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 3);
    regs_read_arr(46)(REG_TRIGGER_OH1_CLUSTER_SIZE_4_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_4_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 4);
    regs_read_arr(47)(REG_TRIGGER_OH1_CLUSTER_SIZE_5_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_5_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 5);
    regs_read_arr(48)(REG_TRIGGER_OH1_CLUSTER_SIZE_6_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_6_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 6);
    regs_read_arr(49)(REG_TRIGGER_OH1_CLUSTER_SIZE_7_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_7_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 7);
    regs_read_arr(50)(REG_TRIGGER_OH1_CLUSTER_SIZE_8_RATE_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_8_RATE_LSB) <= cluster_cnt_rate(1 * 9 + 8);
    regs_read_arr(51)(REG_TRIGGER_OH1_CLUSTER_SIZE_0_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_0_CNT_LSB) <= cluster_cnt(1 * 9 + 0);
    regs_read_arr(52)(REG_TRIGGER_OH1_CLUSTER_SIZE_1_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_1_CNT_LSB) <= cluster_cnt(1 * 9 + 1);
    regs_read_arr(53)(REG_TRIGGER_OH1_CLUSTER_SIZE_2_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_2_CNT_LSB) <= cluster_cnt(1 * 9 + 2);
    regs_read_arr(54)(REG_TRIGGER_OH1_CLUSTER_SIZE_3_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_3_CNT_LSB) <= cluster_cnt(1 * 9 + 3);
    regs_read_arr(55)(REG_TRIGGER_OH1_CLUSTER_SIZE_4_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_4_CNT_LSB) <= cluster_cnt(1 * 9 + 4);
    regs_read_arr(56)(REG_TRIGGER_OH1_CLUSTER_SIZE_5_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_5_CNT_LSB) <= cluster_cnt(1 * 9 + 5);
    regs_read_arr(57)(REG_TRIGGER_OH1_CLUSTER_SIZE_6_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_6_CNT_LSB) <= cluster_cnt(1 * 9 + 6);
    regs_read_arr(58)(REG_TRIGGER_OH1_CLUSTER_SIZE_7_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_7_CNT_LSB) <= cluster_cnt(1 * 9 + 7);
    regs_read_arr(59)(REG_TRIGGER_OH1_CLUSTER_SIZE_8_CNT_MSB downto REG_TRIGGER_OH1_CLUSTER_SIZE_8_CNT_LSB) <= cluster_cnt(1 * 9 + 8);
    regs_read_arr(60)(REG_TRIGGER_OH1_LINK0_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(1)(15 downto 0);
    regs_read_arr(60)(REG_TRIGGER_OH1_LINK1_SBIT_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_SBIT_OVERFLOW_CNT_LSB) <= sbit_overflow_cnt(1)(31 downto 16);
    regs_read_arr(61)(REG_TRIGGER_OH1_LINK0_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH1_LINK0_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(1)(15 downto 0);
    regs_read_arr(61)(REG_TRIGGER_OH1_LINK1_MISSED_COMMA_CNT_MSB downto REG_TRIGGER_OH1_LINK1_MISSED_COMMA_CNT_LSB) <= missed_comma_cnt(1)(31 downto 16);
    regs_read_arr(62)(REG_TRIGGER_OH1_LINK0_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_OVERFLOW_CNT_LSB) <= link_overflow_cnt(1)(15 downto 0);
    regs_read_arr(62)(REG_TRIGGER_OH1_LINK1_OVERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_OVERFLOW_CNT_LSB) <= link_overflow_cnt(1)(31 downto 16);
    regs_read_arr(63)(REG_TRIGGER_OH1_LINK0_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK0_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(1)(15 downto 0);
    regs_read_arr(63)(REG_TRIGGER_OH1_LINK1_UNDERFLOW_CNT_MSB downto REG_TRIGGER_OH1_LINK1_UNDERFLOW_CNT_LSB) <= link_underflow_cnt(1)(31 downto 16);
    regs_read_arr(64)(REG_TRIGGER_OH1_LINK0_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH1_LINK0_SYNC_WORD_CNT_LSB) <= sync_word_cnt(1)(15 downto 0);
    regs_read_arr(64)(REG_TRIGGER_OH1_LINK1_SYNC_WORD_CNT_MSB downto REG_TRIGGER_OH1_LINK1_SYNC_WORD_CNT_LSB) <= sync_word_cnt(1)(31 downto 16);

    -- Connect write signals
    oh_mask <= regs_write_arr(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB);
    sbitmon_link_select <= regs_write_arr(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);
    reset_cnt <= regs_write_pulse_arr(1);
    sbitmon_reset <= regs_write_pulse_arr(5);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(2)(REG_TRIGGER_CTRL_OH_KILL_MASK_MSB downto REG_TRIGGER_CTRL_OH_KILL_MASK_LSB) <= REG_TRIGGER_CTRL_OH_KILL_MASK_DEFAULT;
    regs_defaults(6)(REG_TRIGGER_SBIT_MONITOR_OH_SELECT_MSB downto REG_TRIGGER_SBIT_MONITOR_OH_SELECT_LSB) <= REG_TRIGGER_SBIT_MONITOR_OH_SELECT_DEFAULT;

    -- Define writable regs
    regs_writable_arr(2) <= '1';
    regs_writable_arr(6) <= '1';

    --==== Registers end ============================================================================
        
end trigger_arch;