------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity oh_link_regs is
    generic(
        g_NUM_OF_OHs : integer := 1
    );
    port(
        -- reset
        reset_i                : in  std_logic;
        clk_i                  : in  std_logic;

        -- Link statuses
        oh_link_status_arr_i   : in  t_oh_link_status_arr(g_NUM_OF_OHs - 1 downto 0);

        -- IPbus
        ipb_reset_i            : in  std_logic;
        ipb_clk_i              : in  std_logic;
        ipb_miso_o             : out ipb_rbus;
        ipb_mosi_i             : in  ipb_wbus
    );
end oh_link_regs;

architecture oh_link_regs_arch of oh_link_regs is
    
    --=== resets ===--
    
    signal reset_global         : std_logic;
    signal reset_local          : std_logic;
    signal reset                : std_logic;
    
    --=== counters ===--
    
    signal tk_error_cnt_arr     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal evt_rcvd_cnt_arr     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal sync_tk_tx_ovf_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_tk_tx_unf_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal sync_tk_rx_ovf_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_tk_rx_unf_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
       
    signal sync_tr0_rx_ovf_arr  : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_tr0_rx_unf_arr  : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal sync_tr1_rx_ovf_arr  : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal sync_tr1_rx_unf_arr  : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal tk_not_in_table_arr  : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal tk_disperr_arr       : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal tr0_not_in_table_arr : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal tr0_disperr_arr      : t_std32_array(g_NUM_OF_OHs - 1 downto 0);

    signal tr1_not_in_table_arr : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal tr1_disperr_arr      : t_std32_array(g_NUM_OF_OHs - 1 downto 0);


    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => clk_i,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    i_optohybrids : for i in 0 to g_NUM_OF_OHs - 1 generate

        i_cnt_tk_error : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_error,
                count_o   => tk_error_cnt_arr(i)
            );
    
        i_cnt_evt_rcvd : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).evt_rcvd,
                count_o   => evt_rcvd_cnt_arr(i)
            );    
    
        i_cnt_sync_tk_tx_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_tx_sync_status.ovf,
                count_o   => sync_tk_tx_ovf_arr(i)
            );    
    
        i_cnt_sync_tk_tx_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_tx_sync_status.unf,
                count_o   => sync_tk_tx_unf_arr(i)
            );    
    
        i_cnt_sync_tk_rx_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_rx_sync_status.ovf,
                count_o   => sync_tk_rx_ovf_arr(i)
            );    
    
        i_cnt_sync_tk_rx_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_rx_sync_status.unf,
                count_o   => sync_tk_rx_unf_arr(i)
            );    
    
        i_cnt_sync_tr0_rx_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr0_rx_sync_status.ovf,
                count_o   => sync_tr0_rx_ovf_arr(i)
            );    
    
        i_cnt_sync_tr0_rx_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr0_rx_sync_status.unf,
                count_o   => sync_tr0_rx_unf_arr(i)
            );    
    
        i_cnt_sync_tr1_rx_ovf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr1_rx_sync_status.ovf,
                count_o   => sync_tr1_rx_ovf_arr(i)
            );    
    
        i_cnt_sync_tr1_rx_unf : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr1_rx_sync_status.unf,
                count_o   => sync_tr1_rx_unf_arr(i)
            );    
    
        i_cnt_tk_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_rx_gt_status.not_in_table,
                count_o   => tk_not_in_table_arr(i)
            );
                
        i_cnt_tk_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tk_rx_gt_status.disperr,
                count_o   => tk_disperr_arr(i)
            );
                
        i_cnt_tr0_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr0_rx_gt_status.not_in_table,
                count_o   => tr0_not_in_table_arr(i)
            );
                
        i_cnt_tr0_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr0_rx_gt_status.disperr,
                count_o   => tr0_disperr_arr(i)
            );
                
        i_cnt_tr1_not_in_table : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr1_rx_gt_status.not_in_table,
                count_o   => tr1_not_in_table_arr(i)
            );
                
        i_cnt_tr1_disperr : entity work.counter
            generic map(
                g_COUNTER_WIDTH => 32
            )
            port map(
                ref_clk_i => clk_i,
                reset_i   => reset,
                en_i      => oh_link_status_arr_i(i).tr1_rx_gt_status.disperr,
                count_o   => tr1_disperr_arr(i)
            );
                
    end generate i_optohybrids;
    
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_OH_LINKS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_OH_LINKS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_OH_LINKS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"000";
    regs_addresses(1)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"100";
    regs_addresses(2)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"101";
    regs_addresses(3)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"102";
    regs_addresses(4)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"103";
    regs_addresses(5)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"104";
    regs_addresses(6)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"105";
    regs_addresses(7)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"106";
    regs_addresses(8)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"107";
    regs_addresses(9)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"108";
    regs_addresses(10)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"109";
    regs_addresses(11)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10a";
    regs_addresses(12)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10b";
    regs_addresses(13)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10c";
    regs_addresses(14)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10d";
    regs_addresses(15)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10e";
    regs_addresses(16)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"10f";
    regs_addresses(17)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"200";
    regs_addresses(18)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"201";
    regs_addresses(19)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"202";
    regs_addresses(20)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"203";
    regs_addresses(21)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"204";
    regs_addresses(22)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"205";
    regs_addresses(23)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"206";
    regs_addresses(24)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"207";
    regs_addresses(25)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"208";
    regs_addresses(26)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"209";
    regs_addresses(27)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20a";
    regs_addresses(28)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20b";
    regs_addresses(29)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20c";
    regs_addresses(30)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20d";
    regs_addresses(31)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20e";
    regs_addresses(32)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"20f";
    regs_addresses(33)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"300";
    regs_addresses(34)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"301";
    regs_addresses(35)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"302";
    regs_addresses(36)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"303";
    regs_addresses(37)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"304";
    regs_addresses(38)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"305";
    regs_addresses(39)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"306";
    regs_addresses(40)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"307";
    regs_addresses(41)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"308";
    regs_addresses(42)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"309";
    regs_addresses(43)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30a";
    regs_addresses(44)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30b";
    regs_addresses(45)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30c";
    regs_addresses(46)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30d";
    regs_addresses(47)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30e";
    regs_addresses(48)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"30f";
    regs_addresses(49)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"400";
    regs_addresses(50)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"401";
    regs_addresses(51)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"402";
    regs_addresses(52)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"403";
    regs_addresses(53)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"404";
    regs_addresses(54)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"405";
    regs_addresses(55)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"406";
    regs_addresses(56)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"407";
    regs_addresses(57)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"408";
    regs_addresses(58)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"409";
    regs_addresses(59)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40a";
    regs_addresses(60)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40b";
    regs_addresses(61)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40c";
    regs_addresses(62)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40d";
    regs_addresses(63)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40e";
    regs_addresses(64)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"40f";
    regs_addresses(65)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"500";
    regs_addresses(66)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"501";
    regs_addresses(67)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"502";
    regs_addresses(68)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"503";
    regs_addresses(69)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"504";
    regs_addresses(70)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"505";
    regs_addresses(71)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"506";
    regs_addresses(72)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"507";
    regs_addresses(73)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"508";
    regs_addresses(74)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"509";
    regs_addresses(75)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50a";
    regs_addresses(76)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50b";
    regs_addresses(77)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50c";
    regs_addresses(78)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50d";
    regs_addresses(79)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50e";
    regs_addresses(80)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"50f";
    regs_addresses(81)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"600";
    regs_addresses(82)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"601";
    regs_addresses(83)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"602";
    regs_addresses(84)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"603";
    regs_addresses(85)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"604";
    regs_addresses(86)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"605";
    regs_addresses(87)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"606";
    regs_addresses(88)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"607";
    regs_addresses(89)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"608";
    regs_addresses(90)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"609";
    regs_addresses(91)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60a";
    regs_addresses(92)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60b";
    regs_addresses(93)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60c";
    regs_addresses(94)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60d";
    regs_addresses(95)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60e";
    regs_addresses(96)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"60f";
    regs_addresses(97)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"700";
    regs_addresses(98)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"701";
    regs_addresses(99)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"702";
    regs_addresses(100)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"703";
    regs_addresses(101)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"704";
    regs_addresses(102)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"705";
    regs_addresses(103)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"706";
    regs_addresses(104)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"707";
    regs_addresses(105)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"708";
    regs_addresses(106)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"709";
    regs_addresses(107)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70a";
    regs_addresses(108)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70b";
    regs_addresses(109)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70c";
    regs_addresses(110)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70d";
    regs_addresses(111)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70e";
    regs_addresses(112)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"70f";
    regs_addresses(113)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"800";
    regs_addresses(114)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"801";
    regs_addresses(115)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"802";
    regs_addresses(116)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"803";
    regs_addresses(117)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"804";
    regs_addresses(118)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"805";
    regs_addresses(119)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"806";
    regs_addresses(120)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"807";
    regs_addresses(121)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"808";
    regs_addresses(122)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"809";
    regs_addresses(123)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80a";
    regs_addresses(124)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80b";
    regs_addresses(125)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80c";
    regs_addresses(126)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80d";
    regs_addresses(127)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80e";
    regs_addresses(128)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"80f";
    regs_addresses(129)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"900";
    regs_addresses(130)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"901";
    regs_addresses(131)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"902";
    regs_addresses(132)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"903";
    regs_addresses(133)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"904";
    regs_addresses(134)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"905";
    regs_addresses(135)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"906";
    regs_addresses(136)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"907";
    regs_addresses(137)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"908";
    regs_addresses(138)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"909";
    regs_addresses(139)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90a";
    regs_addresses(140)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90b";
    regs_addresses(141)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90c";
    regs_addresses(142)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90d";
    regs_addresses(143)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90e";
    regs_addresses(144)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"90f";
    regs_addresses(145)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a00";
    regs_addresses(146)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a01";
    regs_addresses(147)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a02";
    regs_addresses(148)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a03";
    regs_addresses(149)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a04";
    regs_addresses(150)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a05";
    regs_addresses(151)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a06";
    regs_addresses(152)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a07";
    regs_addresses(153)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a08";
    regs_addresses(154)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a09";
    regs_addresses(155)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0a";
    regs_addresses(156)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0b";
    regs_addresses(157)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0c";
    regs_addresses(158)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0d";
    regs_addresses(159)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0e";
    regs_addresses(160)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a0f";
    regs_addresses(161)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b00";
    regs_addresses(162)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b01";
    regs_addresses(163)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b02";
    regs_addresses(164)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b03";
    regs_addresses(165)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b04";
    regs_addresses(166)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b05";
    regs_addresses(167)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b06";
    regs_addresses(168)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b07";
    regs_addresses(169)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b08";
    regs_addresses(170)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b09";
    regs_addresses(171)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0a";
    regs_addresses(172)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0b";
    regs_addresses(173)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0c";
    regs_addresses(174)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0d";
    regs_addresses(175)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0e";
    regs_addresses(176)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b0f";
    regs_addresses(177)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c00";
    regs_addresses(178)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c01";
    regs_addresses(179)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c02";
    regs_addresses(180)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c03";
    regs_addresses(181)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c04";
    regs_addresses(182)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c05";
    regs_addresses(183)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c06";
    regs_addresses(184)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c07";
    regs_addresses(185)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c08";
    regs_addresses(186)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c09";
    regs_addresses(187)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0a";
    regs_addresses(188)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0b";
    regs_addresses(189)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0c";
    regs_addresses(190)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0d";
    regs_addresses(191)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0e";
    regs_addresses(192)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c0f";

    -- Connect read signals
    regs_read_arr(1)(REG_OH_LINKS_OH0_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(0);
    regs_read_arr(2)(REG_OH_LINKS_OH0_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH0_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(0);
    regs_read_arr(3)(REG_OH_LINKS_OH0_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(0);
    regs_read_arr(4)(REG_OH_LINKS_OH0_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(0);
    regs_read_arr(5)(REG_OH_LINKS_OH0_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(0);
    regs_read_arr(6)(REG_OH_LINKS_OH0_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(0);
    regs_read_arr(7)(REG_OH_LINKS_OH0_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH0_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(0);
    regs_read_arr(8)(REG_OH_LINKS_OH0_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH0_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(0);
    regs_read_arr(9)(REG_OH_LINKS_OH0_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH0_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(0);
    regs_read_arr(10)(REG_OH_LINKS_OH0_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH0_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(0);
    regs_read_arr(11)(REG_OH_LINKS_OH0_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(0);
    regs_read_arr(12)(REG_OH_LINKS_OH0_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH0_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(0);
    regs_read_arr(13)(REG_OH_LINKS_OH0_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH0_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(0);
    regs_read_arr(14)(REG_OH_LINKS_OH0_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH0_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(0);
    regs_read_arr(15)(REG_OH_LINKS_OH0_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH0_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(0);
    regs_read_arr(16)(REG_OH_LINKS_OH0_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH0_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(0);
    regs_read_arr(17)(REG_OH_LINKS_OH1_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(1);
    regs_read_arr(18)(REG_OH_LINKS_OH1_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH1_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(1);
    regs_read_arr(19)(REG_OH_LINKS_OH1_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(1);
    regs_read_arr(20)(REG_OH_LINKS_OH1_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(1);
    regs_read_arr(21)(REG_OH_LINKS_OH1_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(1);
    regs_read_arr(22)(REG_OH_LINKS_OH1_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(1);
    regs_read_arr(23)(REG_OH_LINKS_OH1_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH1_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(1);
    regs_read_arr(24)(REG_OH_LINKS_OH1_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH1_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(1);
    regs_read_arr(25)(REG_OH_LINKS_OH1_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH1_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(1);
    regs_read_arr(26)(REG_OH_LINKS_OH1_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH1_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(1);
    regs_read_arr(27)(REG_OH_LINKS_OH1_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(1);
    regs_read_arr(28)(REG_OH_LINKS_OH1_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH1_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(1);
    regs_read_arr(29)(REG_OH_LINKS_OH1_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH1_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(1);
    regs_read_arr(30)(REG_OH_LINKS_OH1_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH1_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(1);
    regs_read_arr(31)(REG_OH_LINKS_OH1_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH1_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(1);
    regs_read_arr(32)(REG_OH_LINKS_OH1_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH1_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(1);
    regs_read_arr(33)(REG_OH_LINKS_OH2_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(2);
    regs_read_arr(34)(REG_OH_LINKS_OH2_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH2_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(2);
    regs_read_arr(35)(REG_OH_LINKS_OH2_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(2);
    regs_read_arr(36)(REG_OH_LINKS_OH2_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(2);
    regs_read_arr(37)(REG_OH_LINKS_OH2_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(2);
    regs_read_arr(38)(REG_OH_LINKS_OH2_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(2);
    regs_read_arr(39)(REG_OH_LINKS_OH2_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH2_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(2);
    regs_read_arr(40)(REG_OH_LINKS_OH2_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH2_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(2);
    regs_read_arr(41)(REG_OH_LINKS_OH2_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH2_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(2);
    regs_read_arr(42)(REG_OH_LINKS_OH2_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH2_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(2);
    regs_read_arr(43)(REG_OH_LINKS_OH2_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(2);
    regs_read_arr(44)(REG_OH_LINKS_OH2_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH2_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(2);
    regs_read_arr(45)(REG_OH_LINKS_OH2_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH2_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(2);
    regs_read_arr(46)(REG_OH_LINKS_OH2_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH2_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(2);
    regs_read_arr(47)(REG_OH_LINKS_OH2_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH2_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(2);
    regs_read_arr(48)(REG_OH_LINKS_OH2_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH2_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(2);
    regs_read_arr(49)(REG_OH_LINKS_OH3_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(3);
    regs_read_arr(50)(REG_OH_LINKS_OH3_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH3_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(3);
    regs_read_arr(51)(REG_OH_LINKS_OH3_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(3);
    regs_read_arr(52)(REG_OH_LINKS_OH3_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(3);
    regs_read_arr(53)(REG_OH_LINKS_OH3_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(3);
    regs_read_arr(54)(REG_OH_LINKS_OH3_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(3);
    regs_read_arr(55)(REG_OH_LINKS_OH3_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH3_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(3);
    regs_read_arr(56)(REG_OH_LINKS_OH3_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH3_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(3);
    regs_read_arr(57)(REG_OH_LINKS_OH3_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH3_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(3);
    regs_read_arr(58)(REG_OH_LINKS_OH3_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH3_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(3);
    regs_read_arr(59)(REG_OH_LINKS_OH3_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(3);
    regs_read_arr(60)(REG_OH_LINKS_OH3_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH3_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(3);
    regs_read_arr(61)(REG_OH_LINKS_OH3_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH3_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(3);
    regs_read_arr(62)(REG_OH_LINKS_OH3_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH3_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(3);
    regs_read_arr(63)(REG_OH_LINKS_OH3_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH3_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(3);
    regs_read_arr(64)(REG_OH_LINKS_OH3_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH3_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(3);
    regs_read_arr(65)(REG_OH_LINKS_OH4_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(4);
    regs_read_arr(66)(REG_OH_LINKS_OH4_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH4_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(4);
    regs_read_arr(67)(REG_OH_LINKS_OH4_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(4);
    regs_read_arr(68)(REG_OH_LINKS_OH4_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(4);
    regs_read_arr(69)(REG_OH_LINKS_OH4_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(4);
    regs_read_arr(70)(REG_OH_LINKS_OH4_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(4);
    regs_read_arr(71)(REG_OH_LINKS_OH4_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH4_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(4);
    regs_read_arr(72)(REG_OH_LINKS_OH4_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH4_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(4);
    regs_read_arr(73)(REG_OH_LINKS_OH4_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH4_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(4);
    regs_read_arr(74)(REG_OH_LINKS_OH4_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH4_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(4);
    regs_read_arr(75)(REG_OH_LINKS_OH4_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(4);
    regs_read_arr(76)(REG_OH_LINKS_OH4_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH4_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(4);
    regs_read_arr(77)(REG_OH_LINKS_OH4_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH4_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(4);
    regs_read_arr(78)(REG_OH_LINKS_OH4_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH4_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(4);
    regs_read_arr(79)(REG_OH_LINKS_OH4_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH4_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(4);
    regs_read_arr(80)(REG_OH_LINKS_OH4_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH4_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(4);
    regs_read_arr(81)(REG_OH_LINKS_OH5_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(5);
    regs_read_arr(82)(REG_OH_LINKS_OH5_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH5_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(5);
    regs_read_arr(83)(REG_OH_LINKS_OH5_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(5);
    regs_read_arr(84)(REG_OH_LINKS_OH5_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(5);
    regs_read_arr(85)(REG_OH_LINKS_OH5_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(5);
    regs_read_arr(86)(REG_OH_LINKS_OH5_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(5);
    regs_read_arr(87)(REG_OH_LINKS_OH5_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH5_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(5);
    regs_read_arr(88)(REG_OH_LINKS_OH5_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH5_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(5);
    regs_read_arr(89)(REG_OH_LINKS_OH5_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH5_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(5);
    regs_read_arr(90)(REG_OH_LINKS_OH5_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH5_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(5);
    regs_read_arr(91)(REG_OH_LINKS_OH5_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(5);
    regs_read_arr(92)(REG_OH_LINKS_OH5_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH5_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(5);
    regs_read_arr(93)(REG_OH_LINKS_OH5_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH5_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(5);
    regs_read_arr(94)(REG_OH_LINKS_OH5_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH5_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(5);
    regs_read_arr(95)(REG_OH_LINKS_OH5_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH5_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(5);
    regs_read_arr(96)(REG_OH_LINKS_OH5_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH5_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(5);
    regs_read_arr(97)(REG_OH_LINKS_OH6_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(6);
    regs_read_arr(98)(REG_OH_LINKS_OH6_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH6_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(6);
    regs_read_arr(99)(REG_OH_LINKS_OH6_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(6);
    regs_read_arr(100)(REG_OH_LINKS_OH6_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(6);
    regs_read_arr(101)(REG_OH_LINKS_OH6_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(6);
    regs_read_arr(102)(REG_OH_LINKS_OH6_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(6);
    regs_read_arr(103)(REG_OH_LINKS_OH6_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH6_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(6);
    regs_read_arr(104)(REG_OH_LINKS_OH6_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH6_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(6);
    regs_read_arr(105)(REG_OH_LINKS_OH6_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH6_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(6);
    regs_read_arr(106)(REG_OH_LINKS_OH6_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH6_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(6);
    regs_read_arr(107)(REG_OH_LINKS_OH6_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(6);
    regs_read_arr(108)(REG_OH_LINKS_OH6_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH6_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(6);
    regs_read_arr(109)(REG_OH_LINKS_OH6_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH6_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(6);
    regs_read_arr(110)(REG_OH_LINKS_OH6_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH6_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(6);
    regs_read_arr(111)(REG_OH_LINKS_OH6_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH6_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(6);
    regs_read_arr(112)(REG_OH_LINKS_OH6_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH6_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(6);
    regs_read_arr(113)(REG_OH_LINKS_OH7_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(7);
    regs_read_arr(114)(REG_OH_LINKS_OH7_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH7_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(7);
    regs_read_arr(115)(REG_OH_LINKS_OH7_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(7);
    regs_read_arr(116)(REG_OH_LINKS_OH7_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(7);
    regs_read_arr(117)(REG_OH_LINKS_OH7_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(7);
    regs_read_arr(118)(REG_OH_LINKS_OH7_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(7);
    regs_read_arr(119)(REG_OH_LINKS_OH7_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH7_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(7);
    regs_read_arr(120)(REG_OH_LINKS_OH7_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH7_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(7);
    regs_read_arr(121)(REG_OH_LINKS_OH7_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH7_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(7);
    regs_read_arr(122)(REG_OH_LINKS_OH7_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH7_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(7);
    regs_read_arr(123)(REG_OH_LINKS_OH7_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(7);
    regs_read_arr(124)(REG_OH_LINKS_OH7_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH7_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(7);
    regs_read_arr(125)(REG_OH_LINKS_OH7_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH7_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(7);
    regs_read_arr(126)(REG_OH_LINKS_OH7_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH7_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(7);
    regs_read_arr(127)(REG_OH_LINKS_OH7_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH7_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(7);
    regs_read_arr(128)(REG_OH_LINKS_OH7_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH7_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(7);
    regs_read_arr(129)(REG_OH_LINKS_OH8_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(8);
    regs_read_arr(130)(REG_OH_LINKS_OH8_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH8_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(8);
    regs_read_arr(131)(REG_OH_LINKS_OH8_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(8);
    regs_read_arr(132)(REG_OH_LINKS_OH8_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(8);
    regs_read_arr(133)(REG_OH_LINKS_OH8_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(8);
    regs_read_arr(134)(REG_OH_LINKS_OH8_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(8);
    regs_read_arr(135)(REG_OH_LINKS_OH8_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH8_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(8);
    regs_read_arr(136)(REG_OH_LINKS_OH8_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH8_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(8);
    regs_read_arr(137)(REG_OH_LINKS_OH8_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH8_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(8);
    regs_read_arr(138)(REG_OH_LINKS_OH8_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH8_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(8);
    regs_read_arr(139)(REG_OH_LINKS_OH8_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(8);
    regs_read_arr(140)(REG_OH_LINKS_OH8_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH8_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(8);
    regs_read_arr(141)(REG_OH_LINKS_OH8_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH8_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(8);
    regs_read_arr(142)(REG_OH_LINKS_OH8_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH8_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(8);
    regs_read_arr(143)(REG_OH_LINKS_OH8_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH8_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(8);
    regs_read_arr(144)(REG_OH_LINKS_OH8_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH8_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(8);
    regs_read_arr(145)(REG_OH_LINKS_OH9_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(9);
    regs_read_arr(146)(REG_OH_LINKS_OH9_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH9_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(9);
    regs_read_arr(147)(REG_OH_LINKS_OH9_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(9);
    regs_read_arr(148)(REG_OH_LINKS_OH9_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(9);
    regs_read_arr(149)(REG_OH_LINKS_OH9_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(9);
    regs_read_arr(150)(REG_OH_LINKS_OH9_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(9);
    regs_read_arr(151)(REG_OH_LINKS_OH9_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH9_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(9);
    regs_read_arr(152)(REG_OH_LINKS_OH9_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH9_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(9);
    regs_read_arr(153)(REG_OH_LINKS_OH9_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH9_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(9);
    regs_read_arr(154)(REG_OH_LINKS_OH9_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH9_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(9);
    regs_read_arr(155)(REG_OH_LINKS_OH9_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(9);
    regs_read_arr(156)(REG_OH_LINKS_OH9_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH9_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(9);
    regs_read_arr(157)(REG_OH_LINKS_OH9_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH9_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(9);
    regs_read_arr(158)(REG_OH_LINKS_OH9_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH9_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(9);
    regs_read_arr(159)(REG_OH_LINKS_OH9_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH9_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(9);
    regs_read_arr(160)(REG_OH_LINKS_OH9_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH9_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(9);
    regs_read_arr(161)(REG_OH_LINKS_OH10_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(10);
    regs_read_arr(162)(REG_OH_LINKS_OH10_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH10_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(10);
    regs_read_arr(163)(REG_OH_LINKS_OH10_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(10);
    regs_read_arr(164)(REG_OH_LINKS_OH10_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(10);
    regs_read_arr(165)(REG_OH_LINKS_OH10_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(10);
    regs_read_arr(166)(REG_OH_LINKS_OH10_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(10);
    regs_read_arr(167)(REG_OH_LINKS_OH10_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH10_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(10);
    regs_read_arr(168)(REG_OH_LINKS_OH10_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH10_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(10);
    regs_read_arr(169)(REG_OH_LINKS_OH10_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH10_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(10);
    regs_read_arr(170)(REG_OH_LINKS_OH10_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH10_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(10);
    regs_read_arr(171)(REG_OH_LINKS_OH10_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(10);
    regs_read_arr(172)(REG_OH_LINKS_OH10_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH10_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(10);
    regs_read_arr(173)(REG_OH_LINKS_OH10_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH10_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(10);
    regs_read_arr(174)(REG_OH_LINKS_OH10_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH10_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(10);
    regs_read_arr(175)(REG_OH_LINKS_OH10_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH10_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(10);
    regs_read_arr(176)(REG_OH_LINKS_OH10_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH10_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(10);
    regs_read_arr(177)(REG_OH_LINKS_OH11_TRACK_LINK_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_ERROR_CNT_LSB) <= tk_error_cnt_arr(11);
    regs_read_arr(178)(REG_OH_LINKS_OH11_VFAT_BLOCK_CNT_MSB downto REG_OH_LINKS_OH11_VFAT_BLOCK_CNT_LSB) <= evt_rcvd_cnt_arr(11);
    regs_read_arr(179)(REG_OH_LINKS_OH11_TRACK_LINK_TX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_TX_SYNC_OVF_CNT_LSB) <= sync_tk_tx_ovf_arr(11);
    regs_read_arr(180)(REG_OH_LINKS_OH11_TRACK_LINK_TX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_TX_SYNC_UNF_CNT_LSB) <= sync_tk_tx_unf_arr(11);
    regs_read_arr(181)(REG_OH_LINKS_OH11_TRACK_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tk_rx_ovf_arr(11);
    regs_read_arr(182)(REG_OH_LINKS_OH11_TRACK_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tk_rx_unf_arr(11);
    regs_read_arr(183)(REG_OH_LINKS_OH11_TRIG0_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH11_TRIG0_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr0_rx_ovf_arr(11);
    regs_read_arr(184)(REG_OH_LINKS_OH11_TRIG0_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH11_TRIG0_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr0_rx_unf_arr(11);
    regs_read_arr(185)(REG_OH_LINKS_OH11_TRIG1_LINK_RX_SYNC_OVF_CNT_MSB downto REG_OH_LINKS_OH11_TRIG1_LINK_RX_SYNC_OVF_CNT_LSB) <= sync_tr1_rx_ovf_arr(11);
    regs_read_arr(186)(REG_OH_LINKS_OH11_TRIG1_LINK_RX_SYNC_UNF_CNT_MSB downto REG_OH_LINKS_OH11_TRIG1_LINK_RX_SYNC_UNF_CNT_LSB) <= sync_tr1_rx_unf_arr(11);
    regs_read_arr(187)(REG_OH_LINKS_OH11_TRACK_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_NOT_IN_TABLE_CNT_LSB) <= tk_not_in_table_arr(11);
    regs_read_arr(188)(REG_OH_LINKS_OH11_TRACK_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH11_TRACK_LINK_DISPERR_CNT_LSB) <= tk_disperr_arr(11);
    regs_read_arr(189)(REG_OH_LINKS_OH11_TRIG0_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH11_TRIG0_LINK_NOT_IN_TABLE_CNT_LSB) <= tr0_not_in_table_arr(11);
    regs_read_arr(190)(REG_OH_LINKS_OH11_TRIG0_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH11_TRIG0_LINK_DISPERR_CNT_LSB) <= tr0_disperr_arr(11);
    regs_read_arr(191)(REG_OH_LINKS_OH11_TRIG1_LINK_NOT_IN_TABLE_CNT_MSB downto REG_OH_LINKS_OH11_TRIG1_LINK_NOT_IN_TABLE_CNT_LSB) <= tr1_not_in_table_arr(11);
    regs_read_arr(192)(REG_OH_LINKS_OH11_TRIG1_LINK_DISPERR_CNT_MSB downto REG_OH_LINKS_OH11_TRIG1_LINK_DISPERR_CNT_LSB) <= tr1_disperr_arr(11);

    -- Connect write signals

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults

    -- Define writable regs

    --==== Registers end ============================================================================
    
end oh_link_regs_arch;

