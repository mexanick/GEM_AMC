------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    20:38:00 2016-08-30
-- Module Name:    GEM_TESTS
-- Description:    This module is the entry point for hardware tests e.g. fiber loopback testing with generated data 
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity gem_tests is
    generic(
        g_NUM_GBT_LINKS     : integer
    );
    port(
        -- reset
        reset_i                 : in  std_logic;
        
        -- TTC
        ttc_clk_i               : in  t_ttc_clks;        
        ttc_cmds_i              : in  t_ttc_cmds;
        
        -- Test control
        gbt_loopback_test_en    : in std_logic;
        
        -- GBT links
        gbt_link_ready_i        : in  std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_tx_data_arr_o       : out t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_rx_data_arr_i       : in  t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        
        -- IPbus
        ipb_reset_i             : in  std_logic;
        ipb_clk_i               : in  std_logic;
        ipb_miso_o              : out ipb_rbus;
        ipb_mosi_i              : in  ipb_wbus        
    );
end gem_tests;

architecture Behavioral of gem_tests is

    signal reset_global         : std_logic;
    signal reset_local          : std_logic;
    signal reset                : std_logic;

    signal gbt_loop_sync_done_arr       : std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_mega_word_cnt_arr   : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_error_cnt_arr       : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    ------ Register signals end ----------------------------------------------    

begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --== GBT loopback test ==--
    
    i_gbt_loopback_tests : for i in 0 to g_NUM_GBT_LINKS - 1 generate
    
        i_gbt_loopback_test_single : entity work.gbt_loopback_test
            port map(
                reset_i          => reset or not gbt_loopback_test_en,
                gbt_clk_i        => ttc_clk_i.clk_40,
                gbt_link_ready_i => gbt_link_ready_i(i),
                gbt_tx_data_o    => gbt_tx_data_arr_o(i),
                gbt_rx_data_i    => gbt_rx_data_arr_i(i),
                link_sync_done_o => gbt_loop_sync_done_arr(i),
                mega_word_cnt_o  => gbt_loop_mega_word_cnt_arr(i),
                error_cnt_o      => gbt_loop_error_cnt_arr(i)
            );
    
    end generate;

    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instantiation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_GEM_TESTS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_GEM_TESTS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_GEM_TESTS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults
      );

    -- Addresses
    regs_addresses(0)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0000";
    regs_addresses(1)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0100";
    regs_addresses(2)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0101";
    regs_addresses(3)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0102";
    regs_addresses(4)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0110";
    regs_addresses(5)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0111";
    regs_addresses(6)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0112";
    regs_addresses(7)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0120";
    regs_addresses(8)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0121";
    regs_addresses(9)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0122";
    regs_addresses(10)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0130";
    regs_addresses(11)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0131";
    regs_addresses(12)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0132";
    regs_addresses(13)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0140";
    regs_addresses(14)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0141";
    regs_addresses(15)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0142";
    regs_addresses(16)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0150";
    regs_addresses(17)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0151";
    regs_addresses(18)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0152";
    regs_addresses(19)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0160";
    regs_addresses(20)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0161";
    regs_addresses(21)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0162";
    regs_addresses(22)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0170";
    regs_addresses(23)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0171";
    regs_addresses(24)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0172";
    regs_addresses(25)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0180";
    regs_addresses(26)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0181";
    regs_addresses(27)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0182";
    regs_addresses(28)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0190";
    regs_addresses(29)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0191";
    regs_addresses(30)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0192";
    regs_addresses(31)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01a0";
    regs_addresses(32)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01a1";
    regs_addresses(33)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01a2";
    regs_addresses(34)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01b0";
    regs_addresses(35)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01b1";
    regs_addresses(36)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01b2";
    regs_addresses(37)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01c0";
    regs_addresses(38)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01c1";
    regs_addresses(39)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01c2";
    regs_addresses(40)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01d0";
    regs_addresses(41)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01d1";
    regs_addresses(42)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01d2";
    regs_addresses(43)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01e0";
    regs_addresses(44)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01e1";
    regs_addresses(45)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01e2";
    regs_addresses(46)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01f0";
    regs_addresses(47)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01f1";
    regs_addresses(48)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"01f2";
    regs_addresses(49)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0200";
    regs_addresses(50)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0201";
    regs_addresses(51)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0202";
    regs_addresses(52)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0210";
    regs_addresses(53)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0211";
    regs_addresses(54)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0212";
    regs_addresses(55)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0220";
    regs_addresses(56)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0221";
    regs_addresses(57)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0222";
    regs_addresses(58)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0230";
    regs_addresses(59)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0231";
    regs_addresses(60)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0232";
    regs_addresses(61)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0240";
    regs_addresses(62)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0241";
    regs_addresses(63)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0242";
    regs_addresses(64)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0250";
    regs_addresses(65)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0251";
    regs_addresses(66)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0252";
    regs_addresses(67)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0260";
    regs_addresses(68)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0261";
    regs_addresses(69)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0262";
    regs_addresses(70)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0270";
    regs_addresses(71)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0271";
    regs_addresses(72)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0272";
    regs_addresses(73)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0280";
    regs_addresses(74)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0281";
    regs_addresses(75)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0282";
    regs_addresses(76)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0290";
    regs_addresses(77)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0291";
    regs_addresses(78)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0292";
    regs_addresses(79)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02a0";
    regs_addresses(80)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02a1";
    regs_addresses(81)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02a2";
    regs_addresses(82)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02b0";
    regs_addresses(83)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02b1";
    regs_addresses(84)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02b2";
    regs_addresses(85)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02c0";
    regs_addresses(86)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02c1";
    regs_addresses(87)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02c2";
    regs_addresses(88)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02d0";
    regs_addresses(89)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02d1";
    regs_addresses(90)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02d2";
    regs_addresses(91)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02e0";
    regs_addresses(92)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02e1";
    regs_addresses(93)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02e2";
    regs_addresses(94)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02f0";
    regs_addresses(95)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02f1";
    regs_addresses(96)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"02f2";
    regs_addresses(97)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0300";
    regs_addresses(98)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0301";
    regs_addresses(99)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0302";
    regs_addresses(100)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0310";
    regs_addresses(101)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0311";
    regs_addresses(102)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0312";
    regs_addresses(103)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0320";
    regs_addresses(104)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0321";
    regs_addresses(105)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0322";
    regs_addresses(106)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0330";
    regs_addresses(107)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0331";
    regs_addresses(108)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0332";

    -- Connect read signals
    regs_read_arr(1)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(0);
    regs_read_arr(2)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0);
    regs_read_arr(3)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0);
    regs_read_arr(4)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(1);
    regs_read_arr(5)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1);
    regs_read_arr(6)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1);
    regs_read_arr(7)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(2);
    regs_read_arr(8)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2);
    regs_read_arr(9)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2);
    regs_read_arr(10)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(3);
    regs_read_arr(11)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(3);
    regs_read_arr(12)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(3);
    regs_read_arr(13)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(4);
    regs_read_arr(14)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(4);
    regs_read_arr(15)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(4);
    regs_read_arr(16)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(5);
    regs_read_arr(17)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(5);
    regs_read_arr(18)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(5);
    regs_read_arr(19)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(6);
    regs_read_arr(20)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(6);
    regs_read_arr(21)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(6);
    regs_read_arr(22)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(7);
    regs_read_arr(23)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(7);
    regs_read_arr(24)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(7);
    regs_read_arr(25)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(8);
    regs_read_arr(26)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(8);
    regs_read_arr(27)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(8);
    regs_read_arr(28)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(9);
    regs_read_arr(29)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(9);
    regs_read_arr(30)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(9);
    regs_read_arr(31)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(10);
    regs_read_arr(32)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(10);
    regs_read_arr(33)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(10);
    regs_read_arr(34)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(11);
    regs_read_arr(35)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(11);
    regs_read_arr(36)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(11);
    regs_read_arr(37)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(12);
    regs_read_arr(38)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(12);
    regs_read_arr(39)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(12);
    regs_read_arr(40)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(13);
    regs_read_arr(41)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(13);
    regs_read_arr(42)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(13);
    regs_read_arr(43)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(14);
    regs_read_arr(44)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(14);
    regs_read_arr(45)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(14);
    regs_read_arr(46)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(15);
    regs_read_arr(47)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(15);
    regs_read_arr(48)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(15);
    regs_read_arr(49)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(16);
    regs_read_arr(50)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(16);
    regs_read_arr(51)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(16);
    regs_read_arr(52)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(17);
    regs_read_arr(53)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(17);
    regs_read_arr(54)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(17);
    regs_read_arr(55)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(18);
    regs_read_arr(56)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(18);
    regs_read_arr(57)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(18);
    regs_read_arr(58)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(19);
    regs_read_arr(59)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(19);
    regs_read_arr(60)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(19);
    regs_read_arr(61)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(20);
    regs_read_arr(62)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(20);
    regs_read_arr(63)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(20);
    regs_read_arr(64)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(21);
    regs_read_arr(65)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(21);
    regs_read_arr(66)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(21);
    regs_read_arr(67)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(22);
    regs_read_arr(68)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(22);
    regs_read_arr(69)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(22);
    regs_read_arr(70)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(23);
    regs_read_arr(71)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(23);
    regs_read_arr(72)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(23);
    regs_read_arr(73)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(24);
    regs_read_arr(74)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(24);
    regs_read_arr(75)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(24);
    regs_read_arr(76)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(25);
    regs_read_arr(77)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(25);
    regs_read_arr(78)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(25);
    regs_read_arr(79)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(26);
    regs_read_arr(80)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(26);
    regs_read_arr(81)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(26);
    regs_read_arr(82)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(27);
    regs_read_arr(83)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(27);
    regs_read_arr(84)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(27);
    regs_read_arr(85)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(28);
    regs_read_arr(86)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(28);
    regs_read_arr(87)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(28);
    regs_read_arr(88)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(29);
    regs_read_arr(89)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(29);
    regs_read_arr(90)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(29);
    regs_read_arr(91)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(30);
    regs_read_arr(92)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(30);
    regs_read_arr(93)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(30);
    regs_read_arr(94)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(31);
    regs_read_arr(95)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(31);
    regs_read_arr(96)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(31);
    regs_read_arr(97)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(32);
    regs_read_arr(98)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(32);
    regs_read_arr(99)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(32);
    regs_read_arr(100)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(33);
    regs_read_arr(101)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(33);
    regs_read_arr(102)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(33);
    regs_read_arr(103)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(34);
    regs_read_arr(104)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(34);
    regs_read_arr(105)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(34);
    regs_read_arr(106)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(35);
    regs_read_arr(107)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(35);
    regs_read_arr(108)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(35);

    -- Connect write signals
    -- NOTE: this should be a write pulse (not implemented yet in the generate_registers.py)
    reset_local <= regs_write_arr(0)(REG_GEM_TESTS_CTRL_RESET_BIT);

    -- Defaults

    --==== Registers end ============================================================================

end Behavioral;
