------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    20:38:00 2016-08-30
-- Module Name:    GEM_TESTS
-- Description:    This module is the entry point for hardware tests e.g. fiber loopback testing with generated data 
------------------------------------------------------------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity gem_tests is
    generic(
        g_NUM_GBT_LINKS     : integer;
        g_NUM_OF_OHs        : integer
    );
    port(
        -- reset
        reset_i                     : in  std_logic;
        
        -- TTC
        ttc_clk_i                   : in  t_ttc_clks;        
        ttc_cmds_i                  : in  t_ttc_cmds;
        
        -- Test control
        loopback_gbt_test_en_i      : in std_logic;
        loopback_8b10b_test_en_i    : in std_logic;
        loopback_8b10b_use_trig_i   : in std_logic;
        
        -- 8b10b links
        daq_8b10b_tx_data_arr_o     : out t_gt_8b10b_tx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        daq_8b10b_rx_data_arr_i     : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        trig0_8b10b_rx_data_arr_i   : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        trig1_8b10b_rx_data_arr_i   : in  t_gt_8b10b_rx_data_arr(g_NUM_OF_OHs - 1 downto 0);
        
        -- GBT links
        gbt_link_ready_i            : in  std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_tx_data_arr_o           : out t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        gbt_rx_data_arr_i           : in  t_gbt_frame_array(g_NUM_GBT_LINKS - 1 downto 0);
        
        -- IPbus
        ipb_reset_i                 : in  std_logic;
        ipb_clk_i                   : in  std_logic;
        ipb_miso_o                  : out ipb_rbus;
        ipb_mosi_i                  : in  ipb_wbus        
    );
end gem_tests;

architecture Behavioral of gem_tests is

    -- reset
    signal reset_global                     : std_logic;
    signal reset_local                      : std_logic;
    signal reset                            : std_logic;

    -- control
    signal gbt_loop_through_oh              : std_logic;
    
    -- gbt loopback status
    signal gbt_loop_sync_done_arr           : std_logic_vector(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_mega_word_cnt_arr       : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    signal gbt_loop_error_cnt_arr           : t_std32_array(g_NUM_GBT_LINKS - 1 downto 0);
    
    -- 8b10b status
    signal all_8b10b_loop_mega_word_cnt_arr : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal daq_8b10b_loop_sync_done_arr     : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal daq_8b10b_loop_error_cnt_arr     : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trig0_8b10b_loop_sync_done_arr   : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal trig0_8b10b_loop_error_cnt_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    signal trig1_8b10b_loop_sync_done_arr   : std_logic_vector(g_NUM_OF_OHs - 1 downto 0);
    signal trig1_8b10b_loop_error_cnt_arr   : t_std32_array(g_NUM_OF_OHs - 1 downto 0);
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_GEM_TESTS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------    

begin

    --== Resets ==--
    
    i_reset_sync : entity work.synchronizer
        generic map(
            N_STAGES => 3
        )
        port map(
            async_i => reset_i,
            clk_i   => ttc_clk_i.clk_40,
            sync_o  => reset_global
        );

    reset <= reset_global or reset_local;
    
    --== GBT loopback test ==--
    
    i_gbt_loopback_tests : for i in 0 to g_NUM_GBT_LINKS - 1 generate
    
        i_gbt_loopback_test_single : entity work.gbt_loopback_test
            port map(
                reset_i          => reset or not loopback_gbt_test_en_i,
                gbt_clk_i        => ttc_clk_i.clk_40,
                gbt_link_ready_i => gbt_link_ready_i(i),
                gbt_tx_data_o    => gbt_tx_data_arr_o(i),
                gbt_rx_data_i    => gbt_rx_data_arr_i(i),
                oh_in_the_loop_i => gbt_loop_through_oh,
                link_sync_done_o => gbt_loop_sync_done_arr(i),
                mega_word_cnt_o  => gbt_loop_mega_word_cnt_arr(i),
                error_cnt_o      => gbt_loop_error_cnt_arr(i)
            );
    
    end generate;

    --== 8b10b loopback test ==--
    
    i_8b10b_loopback_tests : for i in 0 to g_NUM_OF_OHs - 1 generate
    
        i_gbt_loopback_test_single : entity work.gt_8b10b_loopback_test
            port map(
                reset_i                 => reset or not loopback_8b10b_test_en_i,
                link_clk_i              => ttc_clk_i.clk_160,
                daq_tx_data_o           => daq_8b10b_tx_data_arr_o(i),
                daq_rx_data_i           => daq_8b10b_rx_data_arr_i(i),
                trig0_rx_data_i         => trig0_8b10b_rx_data_arr_i(i),
                trig1_rx_data_i         => trig1_8b10b_rx_data_arr_i(i),
                use_trig_links          => loopback_8b10b_use_trig_i,
                mega_word_cnt_o         => all_8b10b_loop_mega_word_cnt_arr(i),
                daq_link_sync_done_o    => daq_8b10b_loop_sync_done_arr(i),
                daq_error_cnt_o         => daq_8b10b_loop_error_cnt_arr(i),
                trig0_link_sync_done_o  => trig0_8b10b_loop_sync_done_arr(i),
                trig0_error_cnt_o       => trig0_8b10b_loop_error_cnt_arr(i),
                trig1_link_sync_done_o  => trig1_8b10b_loop_sync_done_arr(i),
                trig1_error_cnt_o       => trig1_8b10b_loop_error_cnt_arr(i)
            );
    
    end generate;
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_GEM_TESTS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_GEM_TESTS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_GEM_TESTS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => ttc_clk_i.clk_40,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"0000";
    regs_addresses(1)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1000";
    regs_addresses(2)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1010";
    regs_addresses(3)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1011";
    regs_addresses(4)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1012";
    regs_addresses(5)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1020";
    regs_addresses(6)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1021";
    regs_addresses(7)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1022";
    regs_addresses(8)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1030";
    regs_addresses(9)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1031";
    regs_addresses(10)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1032";
    regs_addresses(11)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1040";
    regs_addresses(12)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1041";
    regs_addresses(13)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1042";
    regs_addresses(14)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1050";
    regs_addresses(15)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1051";
    regs_addresses(16)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1052";
    regs_addresses(17)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1060";
    regs_addresses(18)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1061";
    regs_addresses(19)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1062";
    regs_addresses(20)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1070";
    regs_addresses(21)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1071";
    regs_addresses(22)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1072";
    regs_addresses(23)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1080";
    regs_addresses(24)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1081";
    regs_addresses(25)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1082";
    regs_addresses(26)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1090";
    regs_addresses(27)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1091";
    regs_addresses(28)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1092";
    regs_addresses(29)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10a0";
    regs_addresses(30)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10a1";
    regs_addresses(31)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10a2";
    regs_addresses(32)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10b0";
    regs_addresses(33)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10b1";
    regs_addresses(34)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10b2";
    regs_addresses(35)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10c0";
    regs_addresses(36)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10c1";
    regs_addresses(37)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10c2";
    regs_addresses(38)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10d0";
    regs_addresses(39)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10d1";
    regs_addresses(40)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10d2";
    regs_addresses(41)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10e0";
    regs_addresses(42)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10e1";
    regs_addresses(43)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10e2";
    regs_addresses(44)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10f0";
    regs_addresses(45)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10f1";
    regs_addresses(46)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"10f2";
    regs_addresses(47)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1100";
    regs_addresses(48)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1101";
    regs_addresses(49)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1102";
    regs_addresses(50)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1110";
    regs_addresses(51)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1111";
    regs_addresses(52)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1112";
    regs_addresses(53)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1120";
    regs_addresses(54)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1121";
    regs_addresses(55)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1122";
    regs_addresses(56)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1130";
    regs_addresses(57)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1131";
    regs_addresses(58)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1132";
    regs_addresses(59)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1140";
    regs_addresses(60)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1141";
    regs_addresses(61)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1142";
    regs_addresses(62)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1150";
    regs_addresses(63)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1151";
    regs_addresses(64)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1152";
    regs_addresses(65)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1160";
    regs_addresses(66)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1161";
    regs_addresses(67)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1162";
    regs_addresses(68)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1170";
    regs_addresses(69)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1171";
    regs_addresses(70)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1172";
    regs_addresses(71)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1180";
    regs_addresses(72)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1181";
    regs_addresses(73)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1182";
    regs_addresses(74)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1190";
    regs_addresses(75)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1191";
    regs_addresses(76)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1192";
    regs_addresses(77)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11a0";
    regs_addresses(78)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11a1";
    regs_addresses(79)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11a2";
    regs_addresses(80)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11b0";
    regs_addresses(81)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11b1";
    regs_addresses(82)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11b2";
    regs_addresses(83)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11c0";
    regs_addresses(84)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11c1";
    regs_addresses(85)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11c2";
    regs_addresses(86)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11d0";
    regs_addresses(87)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11d1";
    regs_addresses(88)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11d2";
    regs_addresses(89)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11e0";
    regs_addresses(90)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11e1";
    regs_addresses(91)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11e2";
    regs_addresses(92)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11f0";
    regs_addresses(93)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11f1";
    regs_addresses(94)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"11f2";
    regs_addresses(95)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1200";
    regs_addresses(96)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1201";
    regs_addresses(97)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1202";
    regs_addresses(98)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1210";
    regs_addresses(99)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1211";
    regs_addresses(100)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1212";
    regs_addresses(101)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1220";
    regs_addresses(102)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1221";
    regs_addresses(103)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1222";
    regs_addresses(104)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1230";
    regs_addresses(105)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1231";
    regs_addresses(106)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1232";
    regs_addresses(107)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1240";
    regs_addresses(108)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1241";
    regs_addresses(109)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"1242";
    regs_addresses(110)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2010";
    regs_addresses(111)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2011";
    regs_addresses(112)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2012";
    regs_addresses(113)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2013";
    regs_addresses(114)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2014";
    regs_addresses(115)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2020";
    regs_addresses(116)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2021";
    regs_addresses(117)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2022";
    regs_addresses(118)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2023";
    regs_addresses(119)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2024";
    regs_addresses(120)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2030";
    regs_addresses(121)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2031";
    regs_addresses(122)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2032";
    regs_addresses(123)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2033";
    regs_addresses(124)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2034";
    regs_addresses(125)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2040";
    regs_addresses(126)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2041";
    regs_addresses(127)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2042";
    regs_addresses(128)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2043";
    regs_addresses(129)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2044";
    regs_addresses(130)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2050";
    regs_addresses(131)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2051";
    regs_addresses(132)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2052";
    regs_addresses(133)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2053";
    regs_addresses(134)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2054";
    regs_addresses(135)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2060";
    regs_addresses(136)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2061";
    regs_addresses(137)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2062";
    regs_addresses(138)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2063";
    regs_addresses(139)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2064";
    regs_addresses(140)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2070";
    regs_addresses(141)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2071";
    regs_addresses(142)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2072";
    regs_addresses(143)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2073";
    regs_addresses(144)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2074";
    regs_addresses(145)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2080";
    regs_addresses(146)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2081";
    regs_addresses(147)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2082";
    regs_addresses(148)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2083";
    regs_addresses(149)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2084";
    regs_addresses(150)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2090";
    regs_addresses(151)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2091";
    regs_addresses(152)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2092";
    regs_addresses(153)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2093";
    regs_addresses(154)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"2094";
    regs_addresses(155)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a0";
    regs_addresses(156)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a1";
    regs_addresses(157)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a2";
    regs_addresses(158)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a3";
    regs_addresses(159)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20a4";
    regs_addresses(160)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b0";
    regs_addresses(161)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b1";
    regs_addresses(162)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b2";
    regs_addresses(163)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b3";
    regs_addresses(164)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20b4";
    regs_addresses(165)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c0";
    regs_addresses(166)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c1";
    regs_addresses(167)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c2";
    regs_addresses(168)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c3";
    regs_addresses(169)(REG_GEM_TESTS_ADDRESS_MSB downto REG_GEM_TESTS_ADDRESS_LSB) <= '0' & x"20c4";

    -- Connect read signals
    regs_read_arr(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT) <= gbt_loop_through_oh;
    regs_read_arr(2)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(0);
    regs_read_arr(3)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(0);
    regs_read_arr(4)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_0_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(0);
    regs_read_arr(5)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(1);
    regs_read_arr(6)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(1);
    regs_read_arr(7)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_1_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(1);
    regs_read_arr(8)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(2);
    regs_read_arr(9)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(2);
    regs_read_arr(10)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_2_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(2);
    regs_read_arr(11)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(3);
    regs_read_arr(12)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(3);
    regs_read_arr(13)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_3_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(3);
    regs_read_arr(14)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(4);
    regs_read_arr(15)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(4);
    regs_read_arr(16)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_4_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(4);
    regs_read_arr(17)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(5);
    regs_read_arr(18)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(5);
    regs_read_arr(19)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_5_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(5);
    regs_read_arr(20)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(6);
    regs_read_arr(21)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(6);
    regs_read_arr(22)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_6_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(6);
    regs_read_arr(23)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(7);
    regs_read_arr(24)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(7);
    regs_read_arr(25)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_7_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(7);
    regs_read_arr(26)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(8);
    regs_read_arr(27)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(8);
    regs_read_arr(28)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_8_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(8);
    regs_read_arr(29)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(9);
    regs_read_arr(30)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(9);
    regs_read_arr(31)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_9_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(9);
    regs_read_arr(32)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(10);
    regs_read_arr(33)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(10);
    regs_read_arr(34)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_10_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(10);
    regs_read_arr(35)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(11);
    regs_read_arr(36)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(11);
    regs_read_arr(37)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_11_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(11);
    regs_read_arr(38)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(12);
    regs_read_arr(39)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(12);
    regs_read_arr(40)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_12_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(12);
    regs_read_arr(41)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(13);
    regs_read_arr(42)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(13);
    regs_read_arr(43)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_13_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(13);
    regs_read_arr(44)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(14);
    regs_read_arr(45)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(14);
    regs_read_arr(46)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_14_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(14);
    regs_read_arr(47)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(15);
    regs_read_arr(48)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(15);
    regs_read_arr(49)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_15_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(15);
    regs_read_arr(50)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(16);
    regs_read_arr(51)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(16);
    regs_read_arr(52)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_16_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(16);
    regs_read_arr(53)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(17);
    regs_read_arr(54)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(17);
    regs_read_arr(55)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_17_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(17);
    regs_read_arr(56)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(18);
    regs_read_arr(57)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(18);
    regs_read_arr(58)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_18_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(18);
    regs_read_arr(59)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(19);
    regs_read_arr(60)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(19);
    regs_read_arr(61)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_19_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(19);
    regs_read_arr(62)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(20);
    regs_read_arr(63)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(20);
    regs_read_arr(64)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_20_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(20);
    regs_read_arr(65)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(21);
    regs_read_arr(66)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(21);
    regs_read_arr(67)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_21_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(21);
    regs_read_arr(68)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(22);
    regs_read_arr(69)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(22);
    regs_read_arr(70)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_22_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(22);
    regs_read_arr(71)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(23);
    regs_read_arr(72)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(23);
    regs_read_arr(73)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_23_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(23);
    regs_read_arr(74)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(24);
    regs_read_arr(75)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(24);
    regs_read_arr(76)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_24_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(24);
    regs_read_arr(77)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(25);
    regs_read_arr(78)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(25);
    regs_read_arr(79)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_25_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(25);
    regs_read_arr(80)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(26);
    regs_read_arr(81)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(26);
    regs_read_arr(82)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_26_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(26);
    regs_read_arr(83)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(27);
    regs_read_arr(84)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(27);
    regs_read_arr(85)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_27_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(27);
    regs_read_arr(86)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(28);
    regs_read_arr(87)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(28);
    regs_read_arr(88)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_28_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(28);
    regs_read_arr(89)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(29);
    regs_read_arr(90)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(29);
    regs_read_arr(91)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_29_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(29);
    regs_read_arr(92)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(30);
    regs_read_arr(93)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(30);
    regs_read_arr(94)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_30_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(30);
    regs_read_arr(95)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(31);
    regs_read_arr(96)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(31);
    regs_read_arr(97)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_31_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(31);
    regs_read_arr(98)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(32);
    regs_read_arr(99)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(32);
    regs_read_arr(100)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_32_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(32);
    regs_read_arr(101)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(33);
    regs_read_arr(102)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(33);
    regs_read_arr(103)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_33_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(33);
    regs_read_arr(104)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(34);
    regs_read_arr(105)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(34);
    regs_read_arr(106)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_34_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(34);
    regs_read_arr(107)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_SYNC_DONE_BIT) <= gbt_loop_sync_done_arr(35);
    regs_read_arr(108)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_MEGA_WORD_CNT_LSB) <= gbt_loop_mega_word_cnt_arr(35);
    regs_read_arr(109)(REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_ERROR_CNT_MSB downto REG_GEM_TESTS_GBT_LOOPBACK_LINK_35_ERROR_CNT_LSB) <= gbt_loop_error_cnt_arr(35);
    regs_read_arr(110)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(0);
    regs_read_arr(110)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(0);
    regs_read_arr(110)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(0);
    regs_read_arr(111)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(0);
    regs_read_arr(112)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(113)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(114)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_0_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(0);
    regs_read_arr(115)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(1);
    regs_read_arr(115)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(1);
    regs_read_arr(115)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(1);
    regs_read_arr(116)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(1);
    regs_read_arr(117)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(1);
    regs_read_arr(118)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(1);
    regs_read_arr(119)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_1_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(1);
    regs_read_arr(120)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(2);
    regs_read_arr(120)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(2);
    regs_read_arr(120)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(2);
    regs_read_arr(121)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(2);
    regs_read_arr(122)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(2);
    regs_read_arr(123)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(2);
    regs_read_arr(124)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_2_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(2);
    regs_read_arr(125)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(3);
    regs_read_arr(125)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(3);
    regs_read_arr(125)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(3);
    regs_read_arr(126)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(3);
    regs_read_arr(127)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(3);
    regs_read_arr(128)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(3);
    regs_read_arr(129)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_3_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(3);
    regs_read_arr(130)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(4);
    regs_read_arr(130)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(4);
    regs_read_arr(130)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(4);
    regs_read_arr(131)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(4);
    regs_read_arr(132)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(4);
    regs_read_arr(133)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(4);
    regs_read_arr(134)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_4_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(4);
    regs_read_arr(135)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(5);
    regs_read_arr(135)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(5);
    regs_read_arr(135)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(5);
    regs_read_arr(136)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(5);
    regs_read_arr(137)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(5);
    regs_read_arr(138)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(5);
    regs_read_arr(139)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_5_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(5);
    regs_read_arr(140)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(6);
    regs_read_arr(140)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(6);
    regs_read_arr(140)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(6);
    regs_read_arr(141)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(6);
    regs_read_arr(142)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(6);
    regs_read_arr(143)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(6);
    regs_read_arr(144)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_6_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(6);
    regs_read_arr(145)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(7);
    regs_read_arr(145)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(7);
    regs_read_arr(145)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(7);
    regs_read_arr(146)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(7);
    regs_read_arr(147)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(7);
    regs_read_arr(148)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(7);
    regs_read_arr(149)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_7_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(7);
    regs_read_arr(150)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(8);
    regs_read_arr(150)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(8);
    regs_read_arr(150)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(8);
    regs_read_arr(151)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(8);
    regs_read_arr(152)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(8);
    regs_read_arr(153)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(8);
    regs_read_arr(154)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_8_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(8);
    regs_read_arr(155)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(9);
    regs_read_arr(155)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(9);
    regs_read_arr(155)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(9);
    regs_read_arr(156)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(9);
    regs_read_arr(157)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(9);
    regs_read_arr(158)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(9);
    regs_read_arr(159)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_9_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(9);
    regs_read_arr(160)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(10);
    regs_read_arr(160)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(10);
    regs_read_arr(160)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(10);
    regs_read_arr(161)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(10);
    regs_read_arr(162)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(10);
    regs_read_arr(163)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(10);
    regs_read_arr(164)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_10_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(10);
    regs_read_arr(165)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_DAQ_SYNC_DONE_BIT) <= daq_8b10b_loop_sync_done_arr(11);
    regs_read_arr(165)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG0_SYNC_DONE_BIT) <= trig0_8b10b_loop_sync_done_arr(11);
    regs_read_arr(165)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG1_SYNC_DONE_BIT) <= trig1_8b10b_loop_sync_done_arr(11);
    regs_read_arr(166)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_MEGA_WORD_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_MEGA_WORD_CNT_LSB) <= all_8b10b_loop_mega_word_cnt_arr(11);
    regs_read_arr(167)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_DAQ_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_DAQ_ERROR_CNT_LSB) <= daq_8b10b_loop_error_cnt_arr(11);
    regs_read_arr(168)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG0_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG0_ERROR_CNT_LSB) <= trig0_8b10b_loop_error_cnt_arr(11);
    regs_read_arr(169)(REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG1_ERROR_CNT_MSB downto REG_GEM_TESTS_8b10b_LOOPBACK_LINK_11_TRIG1_ERROR_CNT_LSB) <= trig1_8b10b_loop_error_cnt_arr(11);

    -- Connect write signals
    gbt_loop_through_oh <= regs_write_arr(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT);

    -- Connect write pulse signals
    reset_local <= regs_write_pulse_arr(0);

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(1)(REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_BIT) <= REG_GEM_TESTS_GBT_LOOPBACK_CTRL_LOOP_THROUGH_OH_DEFAULT;

    -- Define writable regs
    regs_writable_arr(1) <= '1';

    --==== Registers end ============================================================================

end Behavioral;
